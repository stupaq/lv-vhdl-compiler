library ieee;
use ieee.std_logic_1164.all;

entity tiny1 is
    generic (gen1 : integer);
    port (in1 : in std_logic;
        out1 : out std_logic);
end;

architecture behavioral of tiny1 is
begin
end;

